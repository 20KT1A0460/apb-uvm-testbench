`include "sequence_t.sv"
`include "sequence_t_multi_slve_on.sv"
