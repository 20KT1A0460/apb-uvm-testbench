`include "test.sv"
`include "test_error.sv"
`include "test_single_write_read.sv"
`include "test_even_write_read.sv"
`include "test_odd_write_read.sv"
`include "test_full_write_read.sv"
`include "test_multi_slve_on.sv"

