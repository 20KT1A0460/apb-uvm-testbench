 
   `include "../interface/interf.sv"
   `include "../rtl/rtl.v"
  `include "../assertion/ass.sv"

   package uvm_venkatesh_package; 
    `include "uvm_macros.svh"
     import uvm_pkg::*;   
  `include "../seq_item/include.sv"
  `include "../sequence/include.sv"
  `include "../components/include.sv"
  `include "../test/include.sv"
  endpackage
