     `include "sequencer.sv"
     `include "driver.sv"
     `include "imonitor.sv"
     `include "agent1.sv"
     `include "omonitor.sv"
     `include "agent2.sv"
     `include "scoreboard.sv"
     `include "subscriber.sv"
     `include "env.sv"

