`include "seq_item.sv"
`include "seq_item_error.sv"
`include "seq_item_single_write_read.sv"
`include "seq_item_even_write_read.sv"
`include "seq_item_odd_write_read.sv"
`include "seq_item_full_write_read.sv"
`include "seq_item_multi_slve_on.sv"

